/*Copyright 2018-2021 T-Head Semiconductor Co., Ltd.

Licensed under the Apache License, Version 2.0 (the "License");
you may not use this file except in compliance with the License.
You may obtain a copy of the License at

    http://www.apache.org/licenses/LICENSE-2.0

Unless required by applicable law or agreed to in writing, software
distributed under the License is distributed on an "AS IS" BASIS,
WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
See the License for the specific language governing permissions and
limitations under the License.
*/

// &ModuleBeg; @23
module cr_coretim_top_dummy(
  iu_yy_xx_dbgon
);

// &Ports; @24
input        iu_yy_xx_dbgon; 

// &Regs; @25

// &Wires; @26



// //&Force("input", "pad_ctim_refclk"); @29
// &Force("input", "iu_yy_xx_dbgon"); @30
// //&Force("output", "ctim_pad_int_vld"); @31

// &ModuleEnd; @33
endmodule


